<svg xmlns="http://www.w3.org/2000/svg" viewBox="0 0 27 27" height="27" width="27"><title>bear-canister-rentals-white-22.svg</title><rect fill="none" x="0" y="0" width="27" height="27"></rect><rect x="0" y="0" width="27" height="27" rx="4" ry="4" fill="#231f20"></rect><path fill="#ffffff" transform="translate(2 2)" d="M18.9,6.7c0,0-0.1,2.9-2.7,2.7C16.2,9.4,15.9,7,18.9,6.7z"></path><path fill="#ffffff" transform="translate(2 2)" d="M16.9,10.5c0.3-0.3,0.8-0.5,1.3-0.5c1,0,1.8,0.8,1.8,1.8v0.1l0,0c0,0.4-0.2,0.9-0.5,1.5c0,0-0.5,1-0.9,1.4
	l0,0c-0.2,0.2-0.5,0.3-0.8,0.3c-0.4,0-0.7-0.2-0.9-0.5l0,0c-0.2,0.3-0.5,0.5-0.9,0.5c-0.3,0-0.6-0.1-0.8-0.3l0,0
	c-0.4-0.5-0.9-1.4-0.9-1.4c-0.3-0.6-0.4-1.1-0.5-1.5l0,0v-0.1c0-1,0.8-1.8,1.8-1.8C16.1,10,16.5,10.2,16.9,10.5"></path><path fill="#ffffff" transform="translate(2 2)" d="M9.8,9.9L7.4,8.6c0-0.1,0-0.1,0-0.2c0-0.9-0.7-1.7-1.5-1.9H5.1c0-0.1,0.1-0.3,0.1-0.4c0-0.8-0.7-1.5-1.5-1.5
	S2.2,5.3,2.2,6.1v0.1L0,6.6v10.7l2.8-3.2l5.5-0.7c0.6-0.1,1.1-0.4,1.4-0.9l0.6-1.4c0.1-0.1,0.1-0.2,0.1-0.4
	C10.4,10.4,10.1,10.1,9.8,9.9z"></path><path fill="#ffffff" transform="translate(2 2)" d="M16.5,2c-3,0-5.5,0.7-5.5,1.5v15c0,0.8,2.5,1.5,5.5,1.5s5.5-0.7,5.5-1.5v-15C22,2.7,19.5,2,16.5,2z M12,18.4
	v-14C13,4.7,14.6,5,16.5,5C18.4,5,20,4.7,21,4.4v14c-1,0.4-2.6,0.6-4.5,0.6S13,18.8,12,18.4z"></path></svg>
